module hexa_display(SW,HEX);
	input [3:0] SW;
	output [6:0] HEX;

	zero mod0(
		.a(SW[0]),
		.b(SW[1]),
		.c(SW[2]),
		.d(SW[3]),
		.m(HEX[0])
);	
	one mod1(
		.a(SW[0]),
		.b(SW[1]),
		.c(SW[2]),
		.d(SW[3]),
		.m(HEX[1])
);	
	two mod2(
			.a(SW[0]),
			.b(SW[1]),
			.c(SW[2]),
			.d(SW[3]),
			.m(HEX[2])
);	

	three mod3(
			.a(SW[0]),
			.b(SW[1]),
			.c(SW[2]),
			.d(SW[3]),
			.m(HEX[3])
);	

	four mod4(
			.a(SW[0]),
			.b(SW[1]),
			.c(SW[2]),
			.d(SW[3]),
			.m(HEX[4])
);	

	five mod5(
			.a(SW[0]),
			.b(SW[1]),
			.c(SW[2]),
			.d(SW[3]),
			.m(HEX[5])
);	

	six mod6(
			.a(SW[0]),
			.b(SW[1]),
			.c(SW[2]),
			.d(SW[3]),
			.m(HEX[6])
);	

endmodule


module zero(a,b,c,d,m);
	input a;
	input b;
	input c;
	input d;
	output m;

	assign m = ~((~d & ~c & ~b & a) | (~d & c & ~b & ~a) | (d & c & ~b & a) | (d & ~c & b & a))
endmodule

module one(a,b,c,d,m);
	input a;
	input b;
	input c;
	input d;
	output m;

	assign m = ~((~d & c & ~b & a)|(d & c & ~a)|(d & b & a)|(c & b & ~a))
endmodule

module two(a,b,c,d,m);
	input a;
	input b;
	input c;
	input d;
	output m;

	assign m = ~((d & c & ~b & ~a)|(d & c & b)|(~d & ~c & b & ~a))
endmodule

module three(a,b,c,d,m);
	input a;
	input b;
	input c;
	input d;
	output m;

	assign m = ~((~d & ~c & ~b & a)|(~d & c & ~b & ~a)|(c & b & a)|(d & ~c & b & a))
endmodule


module four(a,b,c,d,m);
	input a;
	input b;
	input c;
	input d;
	output m;

	assign m = ~((~d & a)|(~c & ~b & a)|(~d & c & ~b))
endmodule

module five(a,b,c,d,m);
	input a;
	input b;
	input c;
	input d;
	output m;

	assign m = ~((~d & ~c & b)|(~d & ~c & a)|(~d & b & a)|(d & c & ~b & a))
endmodule

module six(a,b,c,d,m);
	input a;
	input b;
	input c;
	input d;
	output m;

	assign m = ~((~d & ~c & ~b)|(d & c & ~b & ~a)|(~d & c & b & a))
endmodule

